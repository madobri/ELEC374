module ALU (
   wire[31:0] ouput; 
);

   

endmodule
