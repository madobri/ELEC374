module orALU(
	input [31:0] A, //32 bit input 1
	input [31:0] B, // 32 bit input 2
	output [63:0] Result //64 bit result
	
);

	assign Result = A|B;
	
endmodule


