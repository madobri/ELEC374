module divisor (
    input clk, reset,                 	// Clock and reset input
    input signed [31:0] M,       // 32 bit Divisor (will be extended to 33-bit)
    input signed [31:0] Q,       // 32 bit Dividend
    output wire [63:0] Result // Quotient + Remainder output
);

    reg [31:0] Q_reg;         // Register to hold the quotient
    reg signed [32:0] A;      // 33 bit accumulator for remainder
    reg signed [32:0] M_neg, M_Pos; // Modified divisor values
    reg signed [32:0] M_extended;   // 33 bit sign-extended divisor
    integer count; // counter for each iteration

    initial count = 0;  

    always @(posedge clk) begin
		 
			if (~reset) begin
				A = 0;  
				Q_reg = 0; 
				count = 0;
			end
			
	 
        else if (count == 0) begin
            count = 1;
				M_extended = {M[31], M};
				
            // Initialize division registers
            A = 33'b0;    
            Q_reg = Q;     

            // Handle signed division cases correctly
            if (M_extended[32] == 1) begin
                M_neg = M_extended;        
                M_Pos = ~M_extended+1;
            end else begin
                M_neg = ~M_extended+1;       
                M_Pos = M_extended;
            end
        end 
        else if (count > 0 && count < 33) begin  // Increased to 33 cycles
            // Shift Left
            {A, Q_reg} = {A, Q_reg} << 1;
	
            // Subtract M from A by adding negative
            A = A + M_neg; 

            // Check sign and restore if necessary
            if (A[32] == 1) begin  
					 Q_reg[0] = 0;   // Append 0 to quotient
                A = A + M_Pos;  // Restore A if it's negative
            end else begin
                Q_reg[0] = 1;   // Append 1 to quotient
            end

            // Increment count to indicate the clock cycle has completed
            count = count + 1; 

        end
    end
	 assign Result = {A[31:0], Q_reg};
endmodule
