module notALU(
	input [31:0] A, //32 bit input
	output [63:0] Result //64 bit result

); 

	assign Result = ~A; 
	
endmodule
